/*
 * 程序功能：74LS138---3线-8线译码器
 * 输入变量 S1：使能端，高电平有效，S2_，S3_：辅助使能端，低电平有效，A：待译码的数字
 * 输出变量 Y_：译码后结果，低电平有效
 */
module Decoder38_74LS138(S1, S2_, S3_, A, Y_);
  input S1, S2_, S3_;
  input [2:0] A;
  output Y_;
  reg [7:0] Y_;
  always @ (S1, S2_, S3_, A)
  begin
    // 总使能端 S = (S1 & ~(~S2_ | ~S3_))无效时，至全部输出为 1
    if(~(S1 & ~(~S2_ | ~S3_)))
      Y_ = 8'hff;
    else
    begin
      Y_[0] = A[0] | A[1] | A[2];
      Y_[1] = ~A[0] | A[1] | A[2];
      Y_[2] = A[0] | ~A[1] | A[2];
      Y_[3] = ~A[0] | ~A[1] | A[2];
      Y_[4] = A[0] | A[1] | ~A[2];
      Y_[5] = ~A[0] | A[1] | ~A[2];
      Y_[6] = A[0] | ~A[1] |~ A[2];
      Y_[7] = ~A[0] | ~A[1] | ~A[2];
    end
  end
endmodule
