/*
 * 程序使用了缩位运算符以使代码紧凑化，为方便阅读，均已单独标出
 * 程序功能：74LS148--8线-3线编码器
 * 输入与输出均为低电平有效
 * 输入变量 S_：使能端，I_：待编码的数字
 * 输出变量 Y_：编码后结果，Ys_、Yex_：表示电路工作状态
 */
module Encoder83_74LS148(S_, I_, Y_, Ys_, Yex_);
  input S_;
  input [7:0] I_;
  output [2:0] Y_;
  output Ys_, Yex_;
  assign Y_[0] = ~(~S_ & (I_[1] & ~I_[2] & ~I_[4] & ~I_[6] | I_[3] & ~I_[4] & ~I_[6] | I_[5] & ~I_[6] | I_[7]));
  // 使用了缩位或运算 & 和 |
  assign Y_[1] = ~(~S_ & (I_[2] & &(~I_[5:4]) | I_[3] & &(~I_[5:4]) | |I_[7:6]));
  // 使用了缩位或运算 |
  assign Y_[2] = ~(~S_ & |I_[7:4]);
  // 使用了缩位与运算 &
  assign Ys_ = ~(~S_ &  &(~I_));
  // 使用了缩位或运算 |
  assign Yex_ = ~(~S_ & |I_);
endmodule
